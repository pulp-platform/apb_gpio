// Copyright 2015 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License”); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

`define REG_PADDIR      6'b000000 //BASEADDR+0x00
`define REG_PADIN       6'b000001 //BASEADDR+0x04
`define REG_PADOUT      6'b000010 //BASEADDR+0x08
`define REG_INTEN       6'b000011 //BASEADDR+0x0C
`define REG_INTTYPE0    6'b000100 //BASEADDR+0x10
`define REG_INTTYPE1    6'b000101 //BASEADDR+0x14
`define REG_INTSTATUS   6'b000110 //BASEADDR+0x18

`define REG_PADCFG0     6'b001000 //BASEADDR+0x20
`define REG_PADCFG1     6'b001001 //BASEADDR+0x24
`define REG_PADCFG2     6'b001010 //BASEADDR+0x28
`define REG_PADCFG3     6'b001011 //BASEADDR+0x2C
`define REG_PADCFG4     6'b001100 //BASEADDR+0x30
`define REG_PADCFG5     6'b001101 //BASEADDR+0x34
`define REG_PADCFG6     6'b001110 //BASEADDR+0x38
`define REG_PADCFG7     6'b001111 //BASEADDR+0x3C

`define REG_INTSTAT_A   6'b010000 //BASEADDR+0x40
`define REG_INTSTAT_B   6'b010001 //BASEADDR+0x44
`define REG_INTSTAT_C   6'b010010 //BASEADDR+0x48
`define REG_INTSTAT_D   6'b010011 //BASEADDR+0x4C

`define REG_TRIPH_IN       6'b010100 //BASEADDR+0x50
`define REG_TRIPH_OUT      6'b010101 //BASEADDR+0x54
`define REG_TRIPH_INTEN    6'b010110 //BASEADDR+0x58
`define REG_TRIPH_INTTYP0  6'b010111 //BASEADDR+0x5C
`define REG_TRIPH_INTTYP1  6'b011000 //BASEADDR+0x60
`define REG_TRIPH_INTSTAT  6'b011001 //BASEADDR+0x64
`define REG_TRIPH_IST_DCDC 6'b011010 //BASEADDR+0x68
`define REG_TRIPH_IST_WAKE 6'b011011 //BASEADDR+0x6C

// `define BLABLA_REG      6'b011100 //BASEADDR+0x70
// `define BLABLA_REG      6'b011101 //BASEADDR+0x74
// `define BLABLA_REG      6'b011110 //BASEADDR+0x78
// `define BLABLA_REG      6'b011111 //BASEADDR+0x7C

`define REG_TEMP_ADC_0     6'b100000 //BASEADDR+0x80
`define REG_TEMP_ADC_1     6'b100001 //BASEADDR+0x84

// Mask for autmatic removal of unused registers
`define GPIO_TRIPH_OUT 32'h81F80000
`define GPIO_TRIPH_IN  ~`GPIO_TRIPH_OUT

module apb_gpio
#(
  parameter APB_ADDR_WIDTH = 12  //APB slaves are 4KB by default
)
(
  input  logic                      HCLK,
  input  logic                      HRESETn,
  input  logic [APB_ADDR_WIDTH-1:0] PADDR,
  input  logic [31:0]               PWDATA,
  input  logic                      PWRITE,
  input  logic                      PSEL,
  input  logic                      PENABLE,
  output logic [31:0]               PRDATA,
  output logic                      PREADY,
  output logic                      PSLVERR,

  input  logic [31:0]               gpio_in,
  output logic [31:0]               gpio_out,
  output logic [31:0]               gpio_dir,
  output logic [31:0][5:0]          gpio_padcfg,
  output logic [3:0]                interrupt,

  output logic                      ana_rstn_o,
  input  logic [17:0]               dcdc_comp_i,
  input  logic                      biendi_sync_i,
  output logic [5:0]                biendi_gp_o,
  input  logic [1:0]                edwin_eoc_i,
  input  logic [1:0]                edwin_ovflow_i,
  input  logic [1:0]                edwin_err_i,
  output logic [11:0]               triphos_events_o,

  input  logic [1:0]                temp_adc_valid_i,
  input  logic [1:0][31:0]          temp_adc_data_i
);

  logic [31:0] r_triphos_inten, r_triphos_intstat;
  logic [31:0] r_triphos_inttype0, r_triphos_inttype1;
  logic [31:0] r_triphos_in, r_triphos_out;
  logic [31:0] r_triphos_sync0, r_triphos_sync1;
  
  logic [1:0]       r_tempadc_valid;
  logic [1:0]       r_tempadc_sync0, r_tempadc_sync1;
  logic [1:0][31:0] r_tempadc_data;

  logic [31:0] s_triphos_in;
  logic [31:0] s_triphos_rise, s_triphos_fall;
  logic [31:0] s_triphos_int_rise, s_triphos_int_fall;
  logic [31:0] s_triphos_int_lev0, s_triphos_int_lev1;
  logic [31:0] s_triphos_int_all;

  logic [1:0]  s_tempadc_valid_rise;

  assign s_triphos_in   = {1'b0,edwin_err_i,edwin_ovflow_i,edwin_eoc_i,6'b0,biendi_sync_i,dcdc_comp_i};
  assign ana_rstn_o     = r_triphos_out[31];
  assign biendi_gp_o    = r_triphos_out[24:19];

  assign s_tempadc_valid_rise = r_tempadc_sync1 & ~r_tempadc_valid;

  assign s_triphos_rise =  r_triphos_sync1 & ~r_triphos_in;
  assign s_triphos_fall = ~r_triphos_sync1 &  r_triphos_in;

  assign s_triphos_int_rise =  r_triphos_inttype1 & ~r_triphos_inttype0 & s_triphos_rise;
  assign s_triphos_int_fall =  r_triphos_inttype1 &  r_triphos_inttype0 & s_triphos_fall;
  assign s_triphos_int_lev0 = ~r_triphos_inttype1 &  r_triphos_inttype0 & ~r_triphos_in;
  assign s_triphos_int_lev1 = ~r_triphos_inttype1 & ~r_triphos_inttype0 &  r_triphos_in;

  assign s_triphos_int_all  = r_triphos_inten & (s_triphos_int_rise | s_triphos_int_fall | s_triphos_int_lev0 | s_triphos_int_lev1);

  logic [31:0] r_gpio_inten;
  logic [31:0] r_gpio_inttype0;
  logic [31:0] r_gpio_inttype1;
  logic [31:0] r_gpio_out;
  logic [31:0] r_gpio_dir;
  logic [31:0] r_gpio_sync0;
  logic [31:0] r_gpio_sync1;
  logic [31:0] r_gpio_in;
  logic [31:0] s_gpio_rise;
  logic [31:0] s_gpio_fall;
  logic [31:0] s_is_int_rise;
  logic [31:0] s_is_int_fall;
  logic [31:0] s_is_int_lev0;
  logic [31:0] s_is_int_lev1;
  logic [31:0] s_is_int_all;
  logic  [3:0] s_rise_int;

  logic  [5:0] s_apb_addr;

  logic [31:0] r_status;

  assign s_apb_addr = PADDR[7:2];

  assign s_gpio_rise = r_gpio_sync1 & ~r_gpio_in; //foreach input check if rising edge
  assign s_gpio_fall = ~r_gpio_sync1 & r_gpio_in; //foreach input check if falling edge

  assign s_is_int_rise =  r_gpio_inttype1 & ~r_gpio_inttype0 & s_gpio_rise; // inttype 01 rise
  assign s_is_int_fall =  r_gpio_inttype1 &  r_gpio_inttype0 & s_gpio_fall; // inttype 00 fall
  assign s_is_int_lev0 = ~r_gpio_inttype1 &  r_gpio_inttype0 & ~r_gpio_in;  // inttype 10 level 0
  assign s_is_int_lev1 = ~r_gpio_inttype1 & ~r_gpio_inttype0 &  r_gpio_in;  // inttype 11 level 1

  //check if bit if interrupt is enabled and if interrupt specified by inttype occurred
  assign s_is_int_all  = r_gpio_inten & (s_is_int_rise | s_is_int_fall | s_is_int_lev0 | s_is_int_lev1);

  //is any bit enabled and specified interrupt happened?
  assign s_rise_int[0] = |s_is_int_all[7:0];
  assign s_rise_int[1] = |s_is_int_all[15:8];
  assign s_rise_int[2] = |s_is_int_all[23:16];
  assign s_rise_int[3] = |s_is_int_all[31:24];

  // assignment of event outputs
  always_comb begin
    triphos_events_o[0] = r_triphos_intstat[18];
    triphos_events_o[1] = r_triphos_intstat[25] | r_triphos_intstat[27];
    triphos_events_o[2] = r_triphos_intstat[26] | r_triphos_intstat[28];
    triphos_events_o[3] = r_triphos_intstat[29] | r_triphos_intstat[30];

    for (int i=0; i<4; i++)
      interrupt[i] = |r_status[i*8 +: 8];

    for (int i=0; i<6; i++)
      triphos_events_o[4+i] = |r_triphos_intstat[i*3 +: 3];

    triphos_events_o[10] = s_tempadc_valid_rise[0];
    triphos_events_o[11] = s_tempadc_valid_rise[1];
  end

  always_ff @(posedge HCLK, negedge HRESETn) begin
    if(~HRESETn) begin
      r_status          <= '0;
      r_triphos_intstat <= '0;
    end
    else begin
      
      for (int i=0; i<2; i++) begin
        if (s_tempadc_valid_rise[i])
          r_tempadc_data[i] <= temp_adc_data_i[i];
      end

      // latch & clear on byte level
      for (int i=0; i<4; i++) begin
        if (PSEL && PENABLE && !PWRITE && (s_apb_addr == (`REG_INTSTAT_A + i)))
          r_status[i*8 +: 8] <= 8'b0;
        else if ( ~(|r_status[i*8 +: 8]) && s_rise_int[i] )
          r_status[i*8 +: 8] <= s_is_int_all[i*8 +: 8];
      end

      if (PSEL && PENABLE && !PWRITE && (s_apb_addr == `REG_TRIPH_IST_DCDC))
        r_triphos_intstat[17:0] <= '0;
      else if ( ~(|r_triphos_intstat[17:0]) && |s_triphos_int_all[17:0] )
        r_triphos_intstat[17:0] <= s_triphos_int_all[17:0];

      if (PSEL && PENABLE && !PWRITE && (s_apb_addr == `REG_TRIPH_IST_WAKE)) begin
        r_triphos_intstat[18]    <= 1'b0;
        r_triphos_intstat[30:25] <= 6'b0;
      end
      else if ( ~(|{r_triphos_intstat[30:25],r_triphos_intstat[18]}) && |{s_triphos_int_all[30:25],s_triphos_int_all[18]} ) begin
        r_triphos_intstat[18]    <= s_triphos_int_all[18];
        r_triphos_intstat[30:25] <= s_triphos_int_all[30:25];
      end

      // complete clear
      if (PSEL && PENABLE && !PWRITE && (s_apb_addr == `REG_INTSTATUS))
        r_status  <= 32'b0;

      if (PSEL && PENABLE && !PWRITE && (s_apb_addr == `REG_TRIPH_INTSTAT))
        r_triphos_intstat <= 32'b0;

    end
  end

  always_ff @(posedge HCLK, negedge HRESETn) begin
    if(~HRESETn) begin
      r_gpio_sync0    <= '0;
      r_gpio_sync1    <= '0;
      r_gpio_in       <= '0;
      r_triphos_sync0 <= '0;
      r_triphos_sync1 <= '0;
      r_triphos_in    <= '0;
      r_tempadc_sync0 <= '0;
      r_tempadc_sync1 <= '0;
      r_tempadc_valid <= '0;
    end
    else begin
      r_gpio_sync0    <= gpio_in;      //first 2 sync for metastability resolving
      r_gpio_sync1    <= r_gpio_sync0;
      r_gpio_in       <= r_gpio_sync1; //last reg used for edge detection
      r_triphos_sync0 <= s_triphos_in;
      r_triphos_sync1 <= r_triphos_sync0;
      r_triphos_in    <= r_triphos_sync1;
      r_tempadc_sync0 <= temp_adc_valid_i;
      r_tempadc_sync1 <= r_tempadc_sync0;
      r_tempadc_valid <= r_tempadc_sync1;
    end
  end

  always_ff @(posedge HCLK, negedge HRESETn) begin
    if(~HRESETn) begin
      r_gpio_inten    <=  '0;
      r_gpio_inttype0 <=  '0;
      r_gpio_inttype1 <=  '0;
      r_gpio_out      <=  '0;
      r_gpio_dir      <=  '0;

      r_triphos_inten    <= '0;
      r_triphos_inttype0 <= '0;
      r_triphos_inttype1 <= '0;
      r_triphos_out      <= '0;

      for (int i=0;i<32;i++) 
        gpio_padcfg[i] <= '0;
    end
    else begin
      if (PSEL && PENABLE && PWRITE) begin
        case (s_apb_addr)
          `REG_PADDIR:   r_gpio_dir      <= PWDATA;
          `REG_PADOUT:   r_gpio_out      <= PWDATA;
          `REG_INTEN:    r_gpio_inten    <= PWDATA;
          `REG_INTTYPE0: r_gpio_inttype0 <= PWDATA;
          `REG_INTTYPE1: r_gpio_inttype1 <= PWDATA;

          `REG_TRIPH_OUT:     r_triphos_out      <= PWDATA & `GPIO_TRIPH_OUT;
          `REG_TRIPH_INTEN:   r_triphos_inten    <= PWDATA & `GPIO_TRIPH_IN;
          `REG_TRIPH_INTTYP0: r_triphos_inttype0 <= PWDATA & `GPIO_TRIPH_IN;
          `REG_TRIPH_INTTYP1: r_triphos_inttype1 <= PWDATA & `GPIO_TRIPH_IN;

          `REG_PADCFG0:
          begin
            gpio_padcfg[0]  <= PWDATA[4:0];
            gpio_padcfg[1]  <= PWDATA[12:8];
            gpio_padcfg[2]  <= PWDATA[20:16];
            gpio_padcfg[3]  <= PWDATA[28:24];
          end
          `REG_PADCFG1:
          begin
            gpio_padcfg[4]  <= PWDATA[4:0];
            gpio_padcfg[5]  <= PWDATA[12:8];
            gpio_padcfg[6]  <= PWDATA[20:16];
            gpio_padcfg[7]  <= PWDATA[28:24];
          end
          `REG_PADCFG2:
          begin
            gpio_padcfg[8]  <= PWDATA[4:0];
            gpio_padcfg[9]  <= PWDATA[12:8];
            gpio_padcfg[10] <= PWDATA[20:16];
            gpio_padcfg[11] <= PWDATA[28:24];
          end
          `REG_PADCFG3:
          begin
            gpio_padcfg[12] <= PWDATA[4:0];
            gpio_padcfg[13] <= PWDATA[12:8];
            gpio_padcfg[14] <= PWDATA[20:16];
            gpio_padcfg[15] <= PWDATA[28:24];
          end
          `REG_PADCFG4:
          begin
            gpio_padcfg[16] <= PWDATA[4:0];
            gpio_padcfg[17] <= PWDATA[12:8];
            gpio_padcfg[18] <= PWDATA[20:16];
            gpio_padcfg[19] <= PWDATA[28:24];
          end
          `REG_PADCFG5:
          begin
            gpio_padcfg[20] <= PWDATA[4:0];
            gpio_padcfg[21] <= PWDATA[12:8];
            gpio_padcfg[22] <= PWDATA[20:16];
            gpio_padcfg[23] <= PWDATA[28:24];
          end
          `REG_PADCFG6:
          begin
            gpio_padcfg[24] <= PWDATA[4:0];
            gpio_padcfg[25] <= PWDATA[12:8];
            gpio_padcfg[26] <= PWDATA[20:16];
            gpio_padcfg[27] <= PWDATA[28:24];
          end
          `REG_PADCFG7:
          begin
            gpio_padcfg[28]  <= PWDATA[4:0];
            gpio_padcfg[29]  <= PWDATA[12:8];
            gpio_padcfg[30]  <= PWDATA[20:16];
            gpio_padcfg[31]  <= PWDATA[28:24];
          end
        endcase
      end
    end
  end

  always_comb begin
    PRDATA = '0;
    if (PSEL & PENABLE & ~PWRITE) begin
      case (s_apb_addr)
        `REG_PADDIR:    PRDATA = r_gpio_dir;
        `REG_PADIN:     PRDATA = r_gpio_in;
        `REG_PADOUT:    PRDATA = r_gpio_out;
        `REG_INTEN:     PRDATA = r_gpio_inten;
        `REG_INTTYPE0:  PRDATA = r_gpio_inttype0;
        `REG_INTTYPE1:  PRDATA = r_gpio_inttype1;
        `REG_INTSTATUS: PRDATA = r_status;

        `REG_INTSTAT_A: PRDATA[7:0] = r_status[7:0];
        `REG_INTSTAT_B: PRDATA[7:0] = r_status[15:8];
        `REG_INTSTAT_C: PRDATA[7:0] = r_status[23:16];
        `REG_INTSTAT_D: PRDATA[7:0] = r_status[31:24];
  
        `REG_TRIPH_IN:      PRDATA = r_triphos_in;
        `REG_TRIPH_OUT:     PRDATA = r_triphos_out;
        `REG_TRIPH_INTEN:   PRDATA = r_triphos_inten;
        `REG_TRIPH_INTTYP0: PRDATA = r_triphos_inttype0;
        `REG_TRIPH_INTTYP1: PRDATA = r_triphos_inttype1;
        `REG_TRIPH_INTSTAT: PRDATA = r_triphos_intstat;

        `REG_TRIPH_IST_DCDC: PRDATA[17:0] = r_triphos_intstat[17:0];
        `REG_TRIPH_IST_WAKE: PRDATA[6:0]  = {r_triphos_intstat[30:25],r_triphos_intstat[18]};
  
        `REG_TEMP_ADC_0:     PRDATA = r_tempadc_data[0];
        `REG_TEMP_ADC_1:     PRDATA = r_tempadc_data[1];

        `REG_PADCFG0:   PRDATA = {2'b00,gpio_padcfg[3], 2'b00,gpio_padcfg[2], 2'b00,gpio_padcfg[1], 2'b00,gpio_padcfg[0]};
        `REG_PADCFG1:   PRDATA = {2'b00,gpio_padcfg[7], 2'b00,gpio_padcfg[6], 2'b00,gpio_padcfg[5], 2'b00,gpio_padcfg[4]};
        `REG_PADCFG2:   PRDATA = {2'b00,gpio_padcfg[11],2'b00,gpio_padcfg[10],2'b00,gpio_padcfg[9], 2'b00,gpio_padcfg[8]};
        `REG_PADCFG3:   PRDATA = {2'b00,gpio_padcfg[15],2'b00,gpio_padcfg[14],2'b00,gpio_padcfg[13],2'b00,gpio_padcfg[12]};
        `REG_PADCFG4:   PRDATA = {2'b00,gpio_padcfg[19],2'b00,gpio_padcfg[18],2'b00,gpio_padcfg[17],2'b00,gpio_padcfg[16]};
        `REG_PADCFG5:   PRDATA = {2'b00,gpio_padcfg[23],2'b00,gpio_padcfg[22],2'b00,gpio_padcfg[21],2'b00,gpio_padcfg[20]};
        `REG_PADCFG6:   PRDATA = {2'b00,gpio_padcfg[27],2'b00,gpio_padcfg[26],2'b00,gpio_padcfg[25],2'b00,gpio_padcfg[24]};
        `REG_PADCFG7:   PRDATA = {2'b00,gpio_padcfg[31],2'b00,gpio_padcfg[30],2'b00,gpio_padcfg[29],2'b00,gpio_padcfg[28]};
        default:        PRDATA = '0;
      endcase
    end
  end

  assign gpio_out = r_gpio_out;
  assign gpio_dir = r_gpio_dir;

  assign PREADY  = 1'b1;
  assign PSLVERR = 1'b0;

endmodule

